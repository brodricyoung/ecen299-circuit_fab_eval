.SUBCKT NOTSIMULATED 1
.ENDS NOTSIMULATED